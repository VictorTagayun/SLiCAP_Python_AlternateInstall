"ExIdriver"
* Z:\mnt\DATA\Cursussen\Courses\ASMPT\Session-2\SLiCAP\cir\ExIdriver.asc
V1 N001 0 V value=0 dc=0 dcvar=0 noise=0
N1 N002 0 N001 N003
E1 N003 0 N004 N005 {A_d}
I1 N004 N005 I value=0 dc=0 dcvar=0 noise={S_i}
V2 N002 N004 V value=0 dc=0 dcvar=0 noise={S_v}
R1 N002 N005 {R_s}
V3 N005 0 V value=0 dc=0 dcvar=0 noise=0
I2 N002 N005 I value=0 dc=0 dcvar=0 noise={4*k*T/R_s}
.backanno
.end
